library verilog;
use verilog.vl_types.all;
entity MotorTest_vlg_vec_tst is
end MotorTest_vlg_vec_tst;
